1c
2dd
2cc
3ccc
