1a
2aa
3aaa

