1c
2cc
2cc
3ccc
