1a
3aaa
