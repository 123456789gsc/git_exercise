dddd 
ddd
