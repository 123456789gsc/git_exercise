1e
2ee
3eee
4eeee
