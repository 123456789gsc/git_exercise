1e
2ee
