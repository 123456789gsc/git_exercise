1b
2bb
