1
:wq
3aaa

